module top(o, a, b, c);
output o;
input a, b, c;
and g1(o, a, b, c);
endmodule
