
module top(clk, a, b, op, oe, y, parity, overflow, greater, is_eq,
     less);
  input clk, oe;
  input [7:0] a, b;
  input [1:0] op;
  output [7:0] y;
  output parity, overflow, greater, is_eq, less;
  wire clk, oe;
  wire [7:0] a, b;
  wire [1:0] op;
  wire [7:0] y;
  wire parity, overflow, greater, is_eq, less;
  wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7;
  wire n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15;
  wire n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23;
  wire n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31;
  wire n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39;
  wire n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47;
  wire n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55;
  wire n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63;
  wire n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71;
  wire n_72, n_74, n_75, n_77, n_78, n_79, n_80, n_81;
  wire n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89;
  wire n_90, n_91, n_92, n_93, n_95, n_96, n_97, n_98;
  wire n_99, n_100, n_101, n_102, n_103, n_104, n_105, n_106;
  wire n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114;
  wire n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122;
  wire n_123, n_124, n_125, n_126, n_127, n_130, n_132, n_133;
  wire n_285, n_286, n_287, n_366;
  wire w, w0, w1, w2;
  nand g6133(n_133, w0, w2);
  nand g4(w2, w1, n_127);
  not g1 (w1, n_112);
  nand g0 (w0, w, n_112);
  not g (w, n_127);
  and g6135 (n_130, n_125, 1'b1, n_68, n_126);
  wire w3;
  nand g6134 (n_127, w3, n_115);
  or g5 (w3, n_114, n_123);
  and g6138 (n_124, n_125, n_120, n_121, n_123);
  and g6141 (n_122, n_125, n_111, n_120, n_121);
  and g6139 (n_119, n_125, n_108, n_120, n_121);
  and g6137 (n_118, n_125, n_113, n_120, n_121);
  and g6136 (n_117, n_125, n_110, n_120, n_121);
  and g6142 (n_116, n_125, n_107, n_120, n_121);
  nand g6140 (n_115, n_114, n_123);
  and g6149 (n_126, n_120, n_121);
  wire w4, w5, w6, w7;
  nand g6147 (n_132, w5, w7);
  nand g9 (w7, w6, n_113);
  not g8 (w6, n_109);
  nand g7 (w5, w4, n_109);
  not g6 (w4, n_113);
  wire w8, w9, w10, w11;
  nand g6148 (n_112, w9, w11);
  nand g13 (w11, w10, n_110);
  not g12 (w10, n_111);
  nand g11 (w9, w8, n_111);
  not g10 (w8, n_110);
  wire w12, w13;
  nand g6145 (n_123, w12, w13, n_36);
  or g15 (w13, n_104, n_25);
  or g14 (w12, op[1], n_103);
  nand g6151 (n_120, op[0], n_106);
  nand g6150 (n_121, n_10, n_105);
  wire w14, w15, w16, w17;
  nand g6152 (n_109, w15, w17);
  nand g19 (w17, w16, n_107);
  not g18 (w16, n_108);
  nand g17 (w15, w14, n_108);
  not g16 (w14, n_107);
  not g6154 (n_106, n_105);
  wire w18, w19;
  nand g6153 (n_111, w18, w19, n_41);
  or g21 (w19, n_104, n_39);
  or g20 (w18, op[1], n_101);
  wire w20, w21;
  and g6155 (n_105, w20, w21);
  nand g23 (w21, a[6], n_65);
  nand g22 (w20, n_44, n_102);
  wire w22, w23, w24, w25;
  nand g6156 (n_103, w23, w25);
  nand g27 (w25, w24, n_102);
  not g26 (w24, n_66);
  nand g25 (w23, w22, n_66);
  not g24 (w22, n_102);
  wire w26, w27;
  nand g6157 (n_108, w26, w27, n_34);
  or g29 (w27, n_104, n_26);
  or g28 (w26, op[1], n_96);
  wire w28;
  nor g6159 (n_102, w28, n_58);
  and g30 (w28, n_24, n_100);
  wire w29, w30, w31, w32;
  nand g6161 (n_101, w30, w32);
  nand g34 (w32, w31, n_100);
  not g33 (w31, n_59);
  nand g32 (w30, w29, n_59);
  not g31 (w29, n_100);
  wire w33, w34;
  and g6158 (n_99, w33, w34);
  nand g36 (w34, n_31, n_83);
  nand g35 (w33, n_97, n_91);
  and g6160 (n_98, n_88, n_97, n_87, n_93);
  wire w35, w36;
  nand g6162 (n_107, w35, w36, n_32);
  or g38 (w36, n_104, n_20);
  or g37 (w35, op[1], n_86);
  wire w37, w38;
  and g6164 (n_100, w37, w38);
  nand g40 (w38, a[4], n_71);
  nand g39 (w37, n_55, n_95);
  wire w39, w40, w41, w42;
  nand g6166 (n_96, w40, w42);
  nand g44 (w42, w41, n_95);
  not g43 (w41, n_72);
  nand g42 (w40, w39, n_72);
  not g41 (w39, n_95);
  not g6167 (n_93, n_92);
  nand g6163 (n_91, n_90, n_89);
  nand g6168 (n_92, n_90, n_84);
  wire w43, w44;
  nand g6170 (n_113, w43, w44, n_33);
  or g46 (w44, n_104, n_57);
  or g45 (w43, op[1], n_81);
  wire w45;
  nand g6169 (n_89, w45, n_88);
  or g47 (w45, n_82, n_87);
  wire w46;
  nor g6171 (n_95, w46, n_60);
  and g48 (w46, n_28, n_85);
  wire w47, w48, w49, w50;
  nand g6174 (n_86, w48, w50);
  nand g52 (w50, w49, n_85);
  not g51 (w49, n_61);
  nand g50 (w48, w47, n_61);
  not g49 (w47, n_85);
  wire w51, w52;
  nand g6172 (n_110, w51, w52, n_35);
  or g54 (w52, n_104, n_38);
  or g53 (w51, op[1], n_77);
  nor g6173 (n_84, n_82, n_74, n_83, n_79);
  nor g6175 (n_87, n_78, n_47, n_75);
  wire w53, w54, w55, w56;
  nand g6177 (n_81, w54, w56);
  nand g58 (w56, w55, n_70);
  not g57 (w55, n_80);
  nand g56 (w54, w53, n_80);
  not g55 (w53, n_70);
  wire w57, w58;
  and g6176 (n_85, w57, w58);
  nand g60 (w58, a[2], n_69);
  nand g59 (w57, n_51, n_80);
  nor g6179 (n_79, n_56, n_78, n_64);
  wire w59, w60, w61, w62;
  nand g6180 (n_77, w60, w62);
  nand g64 (w62, w61, n_63);
  not g63 (w61, n_21);
  nand g62 (w60, w59, n_21);
  not g61 (w59, n_63);
  wire w63;
  nor g6178 (n_75, w63, n_74);
  and g65 (w63, n_46, n_52);
  wire w64, w65;
  and g6189 (n_72, w64, w65);
  nand g67 (w65, n_53, n_71);
  nand g66 (w64, a[4], n_54);
  wire w66, w67;
  and g6190 (n_70, w66, w67);
  nand g69 (w67, n_49, n_69);
  nand g68 (w66, a[2], n_50);
  and g6192 (n_114, n_67, n_68);
  wire w68, w69;
  and g6191 (n_66, w68, w69);
  nand g71 (w69, n_42, n_65);
  nand g70 (w68, a[6], n_43);
  wire w70;
  nor g6184 (n_64, w70, n_19);
  and g72 (w70, b[0], n_17);
  wire w71;
  nor g6181 (n_80, w71, n_30);
  and g73 (w71, n_62, n_22);
  wire w72;
  nand g6185 (n_63, w72, n_62);
  or g74 (w72, a[1], n_29);
  wire w73;
  nor g6186 (n_61, w73, n_60);
  and g75 (w73, a[3], n_27);
  wire w74;
  nor g6187 (n_59, w74, n_58);
  and g76 (w74, a[5], n_23);
  nor g6206 (n_57, n_56, n_8);
  nand g6193 (n_55, n_53, n_54);
  nand g6188 (n_52, a[0], n_1, n_18, n_45);
  nand g6199 (n_51, n_49, n_50);
  wire w75;
  nor g6200 (n_48, w75, n_6);
  and g77 (w75, n_90, n_47);
  wire w76;
  nand g6201 (n_46, w76, n_45);
  or g78 (w76, n_56, n_37);
  nand g6202 (n_44, n_42, n_43);
  nand g6205 (n_67, n_11, n_40);
  nand g6194 (n_68, n_12, n_9);
  nand g6226 (n_41, b[5], a[5], n_40);
  and g6212 (n_39, n_88, n_90);
  nor g6211 (n_38, n_7, n_37);
  nand g6221 (n_36, b[6], a[6], n_40);
  nand g6222 (n_35, b[1], a[1], n_40);
  nand g6223 (n_34, b[4], a[4], n_40);
  nand g6224 (n_33, b[2], a[2], n_40);
  nand g6225 (n_32, b[3], a[3], n_40);
  and g6216 (n_97, n_14, n_31);
  nor g6203 (n_30, a[1], n_29);
  nand g6196 (n_28, a[3], n_27);
  nor g6208 (n_26, n_47, n_82);
  nor g6207 (n_25, n_15, n_13);
  nand g6204 (n_24, a[5], n_23);
  nor g6195 (n_58, a[5], n_23);
  nand g6198 (n_62, a[1], n_29);
  nor g6197 (n_60, a[3], n_27);
  not g6217 (n_22, n_21);
  nor g6213 (n_20, n_78, n_74);
  nand g6214 (n_19, n_18, n_45);
  nor g6209 (n_17, a[0], n_37);
  not g6220 (n_65, n_43);
  not g6219 (n_69, n_50);
  not g6218 (n_71, n_54);
  or g6215 (n_83, n_15, n_16);
  not g6234 (n_14, n_13);
  wire w77;
  nand g6210 (n_12, w77, n_11);
  or g79 (w77, b[0], a[0]);
  wire w78, w79, w80, w81;
  nand g6231 (n_54, w79, w81);
  nand g83 (w81, w80, n_10);
  not g82 (w80, b[4]);
  nand g81 (w79, w78, b[4]);
  not g80 (w78, n_10);
  wire w82, w83, w84, w85;
  nand g6233 (n_43, w83, w85);
  nand g87 (w85, w84, n_10);
  not g86 (w84, b[6]);
  nand g85 (w83, w82, b[6]);
  not g84 (w82, n_10);
  not g6246 (n_40, n_9);
  not g6244 (n_8, n_45);
  not g6243 (n_7, n_18);
  wire w86;
  nand g6230 (n_21, w86, n_11);
  or g88 (w86, b[0], n_10);
  wire w87, w88, w89, w90;
  nand g6232 (n_50, w88, w90);
  nand g92 (w90, w89, n_10);
  not g91 (w89, b[2]);
  nand g90 (w88, w87, b[2]);
  not g89 (w87, n_10);
  not g6245 (n_88, n_6);
  and g6237 (n_15, b[6], n_42);
  nor g6236 (n_16, a[7], n_4);
  nor g6235 (n_13, b[6], n_42);
  wire w91, w92, w93, w94;
  nand g6228 (n_27, w92, w94);
  nand g96 (w94, w93, b[3]);
  not g95 (w93, op[0]);
  nand g94 (w92, w91, op[0]);
  not g93 (w91, b[3]);
  wire w95, w96, w97, w98;
  nand g6227 (n_23, w96, w98);
  nand g100 (w98, w97, b[5]);
  not g99 (w97, op[0]);
  nand g98 (w96, w95, op[0]);
  not g97 (w95, b[5]);
  nand g6247 (n_18, b[1], n_3);
  nor g6239 (n_56, b[2], n_49);
  nand g6252 (n_45, b[2], n_49);
  nand g6241 (n_90, b[5], n_5);
  nor g6254 (n_6, b[5], n_5);
  nand g6255 (n_9, op[1], n_10);
  nand g6238 (n_31, a[7], n_4);
  nor g6250 (n_78, b[3], n_2);
  nor g6251 (n_74, a[3], n_0);
  and g6253 (n_82, b[4], n_53);
  nor g6248 (n_47, b[4], n_53);
  nor g6240 (n_37, b[1], n_3);
  wire w99, w100, w101, w102;
  nand g6229 (n_29, w100, w102);
  nand g104 (w102, w101, b[1]);
  not g103 (w101, op[0]);
  nand g102 (w100, w99, op[0]);
  not g101 (w99, b[1]);
  nand g6249 (n_11, b[0], a[0]);
  nand g6242 (n_104, op[0], op[1]);
  not g6262 (n_2, a[3]);
  not g6257 (n_1, b[0]);
  not g6265 (n_42, a[6]);
  not g6261 (n_10, op[0]);
  not g6266 (n_125, op[1]);
  not g6263 (n_0, b[3]);
  not g6264 (n_3, a[1]);
  not g6258 (n_5, a[5]);
  not g6256 (n_4, b[7]);
  not g6259 (n_53, a[4]);
  not g6260 (n_49, a[2]);
  assign less = n_287;
  assign greater = n_99;
  assign y[0] = n_130;
  assign is_eq = n_98;
  assign y[3] = n_116;
  assign y[5] = n_122;
  assign y[6] = n_124;
  assign y[4] = n_119;
  assign y[1] = n_117;
  assign y[2] = n_118;
  assign parity = n_285;
  assign overflow = n_366;
  assign y[7] = n_366;
  wire w103, w104;
  nand g2 (n_285, w103, w104);
  nand g106 (w104, n_132, n_133);
  or g105 (w103, n_132, n_133);
  not g3 (n_287, n_286);
  wire w105, w106;
  nand g6383 (n_286, w105, w106, n_92);
  or g108 (w106, n_16, n_97);
  or g107 (w105, n_83, n_48);
  and g6462 (n_366, n_125, n_126);
endmodule

