module top(internal_n1, n1)
