module top(o, a, b, c, d,e,f,g,h,i,j,k,l,m,n,p,q,r,s,t,u,v,w,x,y,z,_a,_b,_c,_d,_e,_f,_g,_h,_i,_j,_k,_l);
output o;
input a, b, c, d,e,f,g,h,i,j,k,l,m,n,p,q,r,s,t,u,v,w,x,y,z,_a,_b,_c,_d,_e,_f,_g,_h,_i,_j,_k,_l;
wire n1,n2,n3,n4,n5,n6,n7,n8,n9,n10,n11,n12,n13,n14,n15,n16,n17,n18,n19,n20,n21,n22,n23;
wire n24,n25,n26,n27,n28,n29,n30,n31,n32,n33,n34,n35,n36;
or  g1(n1, a, b);
xor g2(n4, e, f);
and g3(n5, n2, n3);
and g4(n8, n5, n6);
xor g5(n10, n6, n12);
and g6(n9, n10, n11);
and g7(n15, n8, n9);
and g8(o, n15, n16);
and g9(n16, n33, n18);
and g10(n18, n23, n24);
xor g11(n24, n26, n27);
and g12(n7, h, i);
and g13(n14, j, k);
and g14(n13, n14, l);
and g15(n21, _h, n22);
or  g16(n22, p, q);
and g17(n20, t, u);
or  g18(n19, s, n20);
xor g19(n25, w, n28);
xor g20(n28, x, y);
xor g21(n29, z ,n30);
and g22(n30, _a, _b);
or  g23(n31, _e, n32);
or  g24(n32, _f, _g);
and g25(n33, n34, n17);
or  g26(n34, n35, n36);
xor g27(n35, _i, _j);
xor g28(n36, _k, _l);
and M1(n2, n1, c);
and M2(n3, d, n4);
and M3(n6, g, n7);
and M4(n12, n13, m);
and M5(n11, n, n21);
and M6(n17, r, n19);
and M7(n27, _d, n31);
and r1(n23, v, n25);
and r2(n26, n29, _c);
endmodule