module top(o, a, b, c, d, e, f, g, h, i, j, k, l, m, n, p, q, r, s, t, u, v, w, x, y, z, _a, _b, _c, _d, _e, _f, _g, _h,_i,_j,_k,_l);
output o;
input a, b, c, d, e, f, g, h, i, j, k, l, m, n, p, q, r, s, t, u, v, w, x, y, z, _a, _b, _c, _d, _e, _f, _g, _h,_i,_j,_k,_l;
wire n1,n2,n3,n4,n5,n6,n7,n8,n9,n10,n11,n12,n13,n14,n15,n16,n17,n18,n19,n20,n21,n22,n23;
wire n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35;

or  g1(n1, a, b);
or  g2(n3, n2, n4);
and g3(n4, n5, n6);
and g4(n8, n3, n7);
xor g5(n27, e, f);
and g6(n30, _h, n31);
and g7(n28, n29, l);
and g8(n29, j, k);
or  g9(n31, p, q);
and g10(n10, n8, n32);
and g11(n26, h, i);
and g12(o, n10, n11);
and g13(n11, n34, n13);
and g14(n13, n14, n15);
and g15(n14, n16, n17);
or  g16(n24, s, n25);
and g17(n25, u, t);
xor g18(n22, _c, n23);
or  g19(n23, v, w);
or  g20(n21, z, n20);
xor g21(n20, _a, _b);
or  g22(n18, _e, n19);
or  g23(n19, _g, _f);
and g24(n32, n33, n9);
xor g25(n33, _i, _j);
and g26(n34, n35, n12);
xor g27(n35, _k, _l);
and M1(n2, n1, c);
and M2(n7, d, n27);
and M3(n9, g, n26);
and M4(n6, n28, m);
and M5(n5, n, n30);
and M6(n12, r, n24);
and M7(n15, _d, n18);
and g_1(n16, n22, x);
and g_2(n17, y, n21);
endmodule